module half_adder (
input wire a,
input wire b,
input wire c,
output wire sum,
output wire carry );

assign sum = a^b;
assign carry = a&b;
endmodule